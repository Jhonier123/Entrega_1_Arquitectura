----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:46:17 09/26/2017 
-- Design Name: 
-- Module Name:    Instruction_memory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity Instruction_memory is
    Port ( addressim : in  STD_LOGIC_VECTOR (31 downto 0);
           reset : in  STD_LOGIC;
           instruction : out  STD_LOGIC_VECTOR (31 downto 0));
end Instruction_memory;

architecture Behavioral of Instruction_memory is

	type rom_type is array(63 downto 0) of STD_LOGIC_VECTOR (31 downto 0);	

	signal arrayinstructions : rom_type := (
                                       "10100000000100000010000000001111",
													"10100010000100000010000000010001",
													"10100100000001000010000000010000",
													"10010000001001000100000000010010",
													"10110000000100000010000000000000",
													"10110010000100000010000000001000",
													"10100100000100000010000000001010",
													"10100100000100000010011000100000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100000000100000010000000001111",
													"10100010000100000010000000010001",
													"10100100000001000010000000010000",
													"10010000001001000100000000010010",
													"10110000000100000010000000000000",
													"10110010000100000010000000001000",
													"10100100000100000010000000001010",
													"10100100000100000010011000100000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100000000100000010000000001111",
													"10100010000100000010000000010001",
													"10100100000001000010000000010000",
													"10010000001001000100000000010010",
													"10110000000100000010000000000000",
													"10110010000100000010000000001000",
													"10100100000100000010000000001010",
													"10100100000100000010011000100000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100000000100000010000000001111",
													"10100010000100000010000000010001",
													"10100100000001000010000000010000",
													"10010000001001000100000000010010",
													"10110000000100000010000000000000",
													"10110010000100000010000000001000",
													"10100100000100000010000000001010",
													"10100100000100000010011000100000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000",
													"10100100000100000010000000010000"
);

begin
    
	 process(addressim,reset)
		begin
			if(reset = '1') then
				instruction <= (others=>'0');
			else
				instruction<=arrayinstructions(conv_integer(addressim(5 downto 0)));
			end if;
	 end process;


end Behavioral;

